`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02.02.2024 13:12:02
// Design Name: 
// Module Name: ieee754add
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ieee754add();
reg [31:0]a,b;
reg [2:0]op;
reg clk;
wire [31:0]z;
wire gr,ls,eq;
aluunit dut(clk,op,a,b,z,gr,ls,eq);
initial
 begin
 clk=1;
op=3'b110;

#190
 op=3'b000;
 b=32'b10111111010000000000000000000000;
 a=32'b00111111100000000000000000000000;
//a=32'b11000000100000000000000000000000;
//b=32'b11000000000000000000000000000000;
#20
op=3'b001;
b=32'b10111111010000000000000000000000;
a=32'b10111111100000000000000000000000;
//a=32'b01000010111111100001000000000000;
//b=32'b01000001100001111000000000000000;
#20
op=3'b010;
a=32'b11000001001000000000000000000000;
b=32'b01000000000000000000000000000000;
#20
op=3'b011;
b=32'b01000010111111100001000000000000;
a=32'b01000001100001111000000000000000;
#20
op=3'b100;
b=32'b00111111110000000000000000000000;
a=32'b01000000001000000000000000000000;

#100 $stop;
end
always #10 clk=~clk;
endmodule
